module	projectileBitMap	(	
					output	logic	[0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors_enemy,
					output	logic	[0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors_player
					
 ) ;

 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;   


localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 



assign object_colors_player = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hB6 },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hB6, 8'hB6, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hFB, 8'hDB, 8'hDB, 8'hDB, 8'hDA, 8'hB6, 8'hFF, 8'hDA, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF },
{8'hFF, 8'hB6, 8'hFF, 8'hDA, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF },
{8'hFF, 8'hDA, 8'hFF, 8'hFF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF },
{8'hFF, 8'hDA, 8'hFF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hB6, 8'hFF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hB6, 8'hFF, 8'hB6, 8'h96, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'h96, 8'h76, 8'h76, 8'h96, 8'h96, 8'h96, 8'h96, 8'h97, 8'h96, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hB6, 8'hFF, 8'hFF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hDA, 8'hFF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'h72, 8'h96, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'h97, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h96, 8'h76, 8'hBA, 8'hDB, 8'hFF, 8'hFF, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hDA, 8'hDA, 8'hFF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'hDB, 8'hB6, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h72, 8'h72, 8'hBB, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB6, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h72, 8'h96, 8'h9B, 8'h9B, 8'hBA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'h72, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h97, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h96, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h96, 8'h97, 8'hBB, 8'hBB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};


assign object_colors_enemy = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h75, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'h50, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h50, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB9, 8'h94, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h74, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB9, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h74, 8'h75, 8'h55, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h75, 8'h9A, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h74, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h50, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h50, 8'h9A, 8'hFF, 8'hFF, 8'h75, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h74, 8'h74, 8'h75, 8'h75, 8'h50, 8'h50, 8'h50, 8'h74, 8'h74, 8'h50, 8'h51, 8'h51, 8'h51, 8'h50, 8'h74, 8'h50, 8'h50, 8'h50, 8'h75, 8'h75, 8'h50, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h51, 8'h75, 8'hBA, 8'hDA, 8'hDF, 8'hDA, 8'h95, 8'h51, 8'h74, 8'h50, 8'h51, 8'h50, 8'h51, 8'h50, 8'h55, 8'h9A, 8'hDA, 8'hDF, 8'hDA, 8'h9A, 8'h55, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h51, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h75, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h75, 8'h75, 8'h75, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'hDA, 8'hFF, 8'hFF, 8'hBA, 8'h50, 8'h50, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h92, 8'hB6, 8'hFF, 8'hFF, 8'hDF, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h50, 8'h50, 8'h51, 8'hDF, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h50, 8'hBA, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'hBA, 8'h75, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h75, 8'h75, 8'h75, 8'hFF, 8'hFF, 8'h49, 8'h00, 8'h00, 8'h92, 8'hB6, 8'h00, 8'hB6, 8'hFF, 8'hBA, 8'h50, 8'h51, 8'hDF, 8'hFF, 8'h6D, 8'h24, 8'hDB, 8'h49, 8'h00, 8'h00, 8'h92, 8'hFF, 8'hDF, 8'h75, 8'h75, 8'h50, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h95, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h92, 8'hB6, 8'h00, 8'h6D, 8'hFF, 8'hDA, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'h24, 8'h24, 8'hDA, 8'h49, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'h75, 8'h74, 8'h50, 8'h96 },
{8'hFF, 8'hFF, 8'hFF, 8'h95, 8'hFF, 8'hDB, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hDA, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'hFF, 8'hFF, 8'h75, 8'hFF, 8'h9A, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h75, 8'hFF, 8'hFF, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB6, 8'hFF, 8'hBA, 8'h50, 8'h51, 8'hDF, 8'hFF, 8'h6D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hDB, 8'h51, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h51, 8'hDA, 8'hFF, 8'hB6, 8'h24, 8'h00, 8'h00, 8'h00, 8'h6D, 8'hFF, 8'hFF, 8'h75, 8'h74, 8'h74, 8'h96, 8'hFF, 8'hDB, 8'h25, 8'h00, 8'h00, 8'h00, 8'h49, 8'hFF, 8'hFF, 8'h96, 8'h50, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h50, 8'h95, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hDB, 8'h92, 8'h6D, 8'hB6, 8'hFF, 8'hFF, 8'h9A, 8'h50, 8'h94, 8'h94, 8'h51, 8'hDA, 8'hFF, 8'hFF, 8'h92, 8'h6D, 8'h92, 8'hFF, 8'hFF, 8'hDA, 8'h51, 8'h50, 8'hFF, 8'h95, 8'h96 },
{8'hFF, 8'h50, 8'hB9, 8'h50, 8'h50, 8'h75, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h50, 8'h94, 8'h94, 8'h94, 8'h74, 8'h51, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h51, 8'h50, 8'h50, 8'h94, 8'h50, 8'h75 },
{8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h75, 8'h51, 8'h50, 8'h75, 8'hBA, 8'hBA, 8'h96, 8'h75, 8'h50, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h74, 8'h50, 8'h75, 8'h9A, 8'hBA, 8'h9A, 8'h75, 8'h50, 8'h51, 8'h75, 8'hBA, 8'hFF, 8'h75, 8'h96 },
{8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'hBA, 8'hDA, 8'hBA, 8'h95, 8'h75, 8'h75, 8'h75, 8'h75, 8'h74, 8'h74, 8'h50, 8'h94, 8'h94, 8'h94, 8'h94, 8'h74, 8'h75, 8'h75, 8'h75, 8'h55, 8'h95, 8'hBA, 8'hDA, 8'hBA, 8'h96, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h51, 8'h95, 8'hDA, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDE, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hBA, 8'h95, 8'h55, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'h75, 8'h95, 8'h75, 8'h50, 8'h50, 8'h50, 8'h50, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h50, 8'h50, 8'h50, 8'h50, 8'h75, 8'h95, 8'h50, 8'hFF },
{8'hFF, 8'h51, 8'h74, 8'h95, 8'h51, 8'h50, 8'h51, 8'h50, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h50, 8'h50, 8'h50, 8'h51, 8'h95, 8'h74, 8'h50, 8'hFF },
{8'hFF, 8'h9A, 8'h50, 8'hFF, 8'h95, 8'h50, 8'h51, 8'h50, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h50, 8'h50, 8'h50, 8'h75, 8'hFF, 8'h75, 8'h75, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h51, 8'h50, 8'h50, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h50, 8'h74, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h74, 8'h50, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h50, 8'h74, 8'h94, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h51, 8'h74, 8'h95, 8'hBA, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h96, 8'h75, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h50, 8'hBA, 8'hDA, 8'h75, 8'h95, 8'hBA, 8'hBA, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDA, 8'hBA, 8'hBA, 8'h95, 8'h75, 8'hBA, 8'hFF, 8'h75, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h50, 8'h74, 8'h94, 8'h51, 8'h75, 8'h51, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h74, 8'h75, 8'h50, 8'h50, 8'h50, 8'h50, 8'h74, 8'h50, 8'h50, 8'h50, 8'h51, 8'h74, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h50, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h75, 8'h94, 8'h95, 8'h9A, 8'hFF, 8'hBA, 8'h74, 8'h50, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h95, 8'hFF, 8'hFF, 8'h75, 8'h50, 8'h50, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h51, 8'h50, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};

endmodule